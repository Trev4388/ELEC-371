library verilog;
use verilog.vl_types.all;
entity processor_vlg_vec_tst is
end processor_vlg_vec_tst;
